// SPDX-License-Identifier: MPL-2.0
//
// rv32i.vh -- rv32i base integer instruction set
// Copyright (C) 2025  Jacob Koziej <jacobkoziej@gmail.com>

`ifndef KEEN_INSTRUCTION_SET_RV32I
`define KEEN_INSTRUCTION_SET_RV32I

// verilog_format: off

// 2.4.1. Integer Register-Immediate Instructions
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_OP_IMM 7'b0010011

`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_ADDI  3'b000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SLTI  3'b010
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SLTIU 3'b011
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_XORI  3'b100
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_ORI   3'b110
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_ANDI  3'b111
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SLLI  3'b001
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SRLI  3'b101
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SRAI  3'b101

`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_LUI   7'b0110111
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_AUIPC 7'b0010111

// 2.4.2. Integer Register-Register Operations
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_OP 7'b0110011

`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_ADD  3'b000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SUB  3'b000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SLL  3'b001
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SLT  3'b010
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SLTU 3'b011
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_XOR  3'b100
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SRL  3'b101
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SRA  3'b101
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_OR   3'b110
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_AND  3'b111

`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_ADD  7'b0000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_SUB  7'b0100000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_SLL  7'b0000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_SLT  7'b0000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_SLTU 7'b0000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_XOR  7'b0000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_SRL  7'b0000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_SRA  7'b0100000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_OR   7'b0000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT7_AND  7'b0000000

// 2.5.1. Unconditional Jumps
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_JAL  7'b1101111
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_JALR 7'b1100111

// 2.5.2. Conditional Branches
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_BRANCH 7'b1100011

`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_BEQ  3'b000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_BNE  3'b001
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_BLT  3'b100
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_BGE  3'b101
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_BLTU 3'b110
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_BGEU 3'b111

// 2.6. Load and Store Instructions
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_LOAD  7'b0000011
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_STORE 7'b0100011

`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_LB  3'b000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_LH  3'b001
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_LW  3'b010
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_LBU 3'b100
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_LHU 3'b101
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SB  3'b000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SH  3'b001
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_SW  3'b010

// 2.7. Memory Ordering Instructions
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_MISC_MEM 7'b0001111

`define KEEN_INSTRUCTION_SET_RV32I_FUNCT3_FENCE 3'b000

// 2.8. Environment Call and Breakpoints
`define KEEN_INSTRUCTION_SET_RV32I_OPCODE_SYSTEM 7'b1110011

`define KEEN_INSTRUCTION_SET_RV32I_FUNCT12_ECALL  12'b000000000000
`define KEEN_INSTRUCTION_SET_RV32I_FUNCT12_EBREAK 12'b000000000001

// verilog_format: on

`endif  // KEEN_INSTRUCTION_SET_RV32I
