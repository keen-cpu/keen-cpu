// SPDX-License-Identifier: MPL-2.0
//
// format.vh -- instruction format
// Copyright (C) 2025  Jacob Koziej <jacobkoziej@gmail.com>

`ifndef KEEN_INSTRUCTION_SET_FORMAT
`define KEEN_INSTRUCTION_SET_FORMAT

// common
`define KEEN_INSTRUCTION_SET_FORMAT_OPCODE_LSB 0
`define KEEN_INSTRUCTION_SET_FORMAT_OPCODE_MSB 6
`define KEEN_INSTRUCTION_SET_FORMAT_RD_LSB 7
`define KEEN_INSTRUCTION_SET_FORMAT_RD_MSB 11
`define KEEN_INSTRUCTION_SET_FORMAT_FUNCT3_LSB 12
`define KEEN_INSTRUCTION_SET_FORMAT_FUNCT3_MSB 14
`define KEEN_INSTRUCTION_SET_FORMAT_RS1_LSB 15
`define KEEN_INSTRUCTION_SET_FORMAT_RS1_MSB 19
`define KEEN_INSTRUCTION_SET_FORMAT_RS2_LSB 20
`define KEEN_INSTRUCTION_SET_FORMAT_RS2_MSB 24

// r-type
`define KEEN_INSTRUCTION_SET_FORMAT_R_TYPE_FUNCT7_LSB 25
`define KEEN_INSTRUCTION_SET_FORMAT_R_TYPE_FUNCT7_MSB 31

// i-type
`define KEEN_INSTRUCTION_SET_FORMAT_I_TYPE_IMM_11_0_LSB 20
`define KEEN_INSTRUCTION_SET_FORMAT_I_TYPE_IMM_11_0_MSB 31

// s-type
`define KEEN_INSTRUCTION_SET_FORMAT_S_TYPE_IMM_4_0_LSB 7
`define KEEN_INSTRUCTION_SET_FORMAT_S_TYPE_IMM_4_0_MSB 11
`define KEEN_INSTRUCTION_SET_FORMAT_S_TYPE_IMM_11_5_LSB 25
`define KEEN_INSTRUCTION_SET_FORMAT_S_TYPE_IMM_11_5_MSB 31

// b-type
`define KEEN_INSTRUCTION_SET_FORMAT_B_TYPE_IMM_11_BIT 7
`define KEEN_INSTRUCTION_SET_FORMAT_B_TYPE_IMM_4_1_LSB 8
`define KEEN_INSTRUCTION_SET_FORMAT_B_TYPE_IMM_4_1_MSB 11
`define KEEN_INSTRUCTION_SET_FORMAT_B_TYPE_IMM_10_5_LSB 25
`define KEEN_INSTRUCTION_SET_FORMAT_B_TYPE_IMM_10_5_MSB 30
`define KEEN_INSTRUCTION_SET_FORMAT_B_TYPE_IMM_12_BIT 31

// u-type
`define KEEN_INSTRUCTION_SET_FORMAT_U_TYPE_IMM_31_12_LSB 12
`define KEEN_INSTRUCTION_SET_FORMAT_U_TYPE_IMM_31_12_MSB 31

// j-type
`define KEEN_INSTRUCTION_SET_FORMAT_J_TYPE_IMM_19_12_LSB 12
`define KEEN_INSTRUCTION_SET_FORMAT_J_TYPE_IMM_19_12_MSB 19
`define KEEN_INSTRUCTION_SET_FORMAT_J_TYPE_IMM_11_BIT 20
`define KEEN_INSTRUCTION_SET_FORMAT_J_TYPE_IMM_10_1_LSB 21
`define KEEN_INSTRUCTION_SET_FORMAT_J_TYPE_IMM_10_1_MSB 30
`define KEEN_INSTRUCTION_SET_FORMAT_J_TYPE_IMM_20_BIT 31

`endif  // KEEN_INSTRUCTION_SET_FORMAT
